-- dasda.vhd

-- Generated using ACDS version 13.0sp1 232 at 2019.10.02.21:51:18

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity dasda is
	port (
		clk_clk       : in std_logic := '0'; --   clk.clk
		reset_reset_n : in std_logic := '0'  -- reset.reset_n
	);
end entity dasda;

architecture rtl of dasda is
begin

end architecture rtl; -- of dasda
