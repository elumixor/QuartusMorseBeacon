// dasda.v

// Generated using ACDS version 13.0sp1 232 at 2019.10.02.21:51:20

`timescale 1 ps / 1 ps
module dasda (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

endmodule
